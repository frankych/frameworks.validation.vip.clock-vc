interface sideband_interface;
    bit side_rst_b;
    bit agent_rst_b;
endinterface