`include "base_pmsb_sequence.sv"
`include "reset_flow_control_sequences.sv"
`include "pmsb_svid_sequences.sv"
`include "pmsb_send_power_state_req_seq.sv"
`include "pmsb_reset_go_messages.sv"
`include "pmsb_reg_read_sequence.sv"
`include "pmsb_reg_write_sequence.sv"
`include "pmsb_send_cmp_msg_sequence.sv"
`include "pmsb_send_cmpd_msg_sequence.sv"