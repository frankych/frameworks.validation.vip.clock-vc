
`ifdef INTEL_SIMONLY
  // saola is filtered for Emulation, 
  // but needs to be present for EmulationSimulation
  // import sla_pkg::*;
`endif
